module strTo7seg (
    input [4:0] A,
    output reg [6:0] SEG
);

always @(*) begin
    case(A)
        5'b00000: SEG = 7'b0111111; //0 : 0
        5'b00001: SEG = 7'b0000110; //1 : 1
        5'b00010: SEG = 7'b1011011; //2 : 2
        5'b00011: SEG = 7'b1001111; //3 : 3
        5'b00100: SEG = 7'b1100110; //4 : 4
        5'b00101: SEG = 7'b1101101; //5 : 5
        5'b00110: SEG = 7'b1111101; //6 : 6
        5'b00111: SEG = 7'b0000111; //7 : 7
        5'b01000: SEG = 7'b1111111; //8 : 8
        5'b01001: SEG = 7'b1101111; //9 : 9
        5'b01010: SEG = 7'b1110111; //10 : A
        5'b01011: SEG = 7'b1111100; //11 : B
        5'b01100: SEG = 7'b0111001; //12 : C
        5'b01101: SEG = 7'b1011110; //13 : D
        5'b01110: SEG = 7'b1111001; //14 : E
        5'b01111: SEG = 7'b1110001; //15 : F
        5'b10000: SEG = 7'b0111101; //16 : G
        5'b10001: SEG = 7'b1110110; //17 : H
        5'b10010: SEG = 7'b0011110; //18: J
        5'b10011: SEG = 7'b0111000; //19 : L
        5'b10100: SEG = 7'b0110111; //20 : N
        5'b10101: SEG = 7'b0111111; //21 : 0
        5'b10110: SEG = 7'b1110011; //22 : P
        5'b10111: SEG = 7'b1010000; ///23 : r
        5'b11000: SEG = 7'b0111110; //24 : U
        5'b11001: SEG = 7'b1101101; //25 : S
        5'b11010: SEG = 7'b1101101; //26 : u
        5'b11011: SEG = 7'b0000000; //27 : spacja
        default: SEG = 7'b0000000; //28 : -
    endcase
end
endmodule