--preskaler