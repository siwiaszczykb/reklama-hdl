module prescaler (
    input wire clk,
    output wire clk1Hz
);

always @(*) begin
    
end

endmodule