--rejestr