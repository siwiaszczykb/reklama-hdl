library IEEE;
use IEEE.std_logic_1164.all;

entity reklama is
port (clk: in std_logic;
		display0: in std_logic_vector(5 downto 0);
		display1: in std_logic_vector(5 downto 0);
		display2: in std_logic_vector(5 downto 0);
		display3: in std_logic_vector(5 downto 0);
		display4: in std_logic_vector(5 downto 0);
		display5: in std_logic_vector(5 downto 0) );
end reklama;

architecture scroll of reklama is 

end scroll;