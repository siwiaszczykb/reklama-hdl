module msg (
    input [3:0] A,
    output reg [4:0] Q
);

always @(*) begin
    case(A)
        4'b0001: Q = 5'b10011; //0 : 19/L
        4'b0010: Q = 5'b11000; //1 : 24/U
        4'b0011: Q = 5'b01011; //2 : 11/B
        4'b0100: Q = 5'b10011; //3 : 19/L
        4'b0101: Q = 5'b00001; //4 : 1/I
        4'b0110: Q = 5'b10100; //5 : 20/N
        4'b0111: Q = 5'b00001; //6 : 1/I
        4'b1000: Q = 5'b01110; //7 : 14/E
        4'b1001: Q = 5'b01100; //8 : 12/C
        4'b1010: Q = 5'b11011; //9 : 27/spacja
        4'b1011: Q = 5'b00010; //10 : 2/2
        4'b1100: Q = 5'b00000; //11 : 0/0
        4'b1101: Q = 5'b00010; //12 : 2/2
        4'b1110: Q = 5'b00101; //13 : 5/5
        4'b1111: Q = 5'b11011; //14 : 27/spacja
        default: Q = 5'b11011; //domyslnie : 27/spacja
    endcase
end
endmodule